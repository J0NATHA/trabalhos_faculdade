CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 71 1536 816
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
80 C:\Users\jonat\AppData\Local\Temp\Rar$EXa10028.42639\CIRCUIT MAKER_CM60S\BOM.DAT
0 7
0 71 1536 816
143654930 0
0
6 Title:
5 Name:
0
0
0
24
13 Logic Switch~
5 97 59 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 59 58 0 1 11
0 6
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
9 2-In NOR~
219 250 377 0 3 22
0 6 8 7
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
3618 0 0
0
0
9 Inverter~
13 176 397 0 2 22
0 4 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
6153 0 0
0
0
9 2-In NOR~
219 346 410 0 3 22
0 7 3 2
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
5394 0 0
0
0
9 2-In NOR~
219 243 451 0 3 22
0 5 4 3
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7734 0 0
0
0
9 Inverter~
13 179 445 0 2 22
0 6 5
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
9914 0 0
0
0
14 Logic Display~
6 435 389 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3747 0 0
0
0
14 Logic Display~
6 436 267 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3549 0 0
0
0
9 Inverter~
13 180 323 0 2 22
0 6 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
7931 0 0
0
0
9 2-In NOR~
219 244 329 0 3 22
0 11 4 10
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
9325 0 0
0
0
9 Inverter~
13 396 288 0 2 22
0 13 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
8903 0 0
0
0
9 2-In NOR~
219 347 288 0 3 22
0 12 10 13
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
3834 0 0
0
0
9 Inverter~
13 177 275 0 2 22
0 4 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
3363 0 0
0
0
9 2-In NOR~
219 251 255 0 3 22
0 6 14 12
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
7668 0 0
0
0
9 Inverter~
13 317 166 0 2 22
0 16 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
4718 0 0
0
0
9 2-In NOR~
219 248 183 0 3 22
0 18 17 16
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
3874 0 0
0
0
9 Inverter~
13 192 167 0 2 22
0 6 18
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
6671 0 0
0
0
9 Inverter~
13 201 202 0 2 22
0 4 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
3789 0 0
0
0
14 Logic Display~
6 362 146 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4871 0 0
0
0
14 Logic Display~
6 277 74 0 1 2
10 19
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3750 0 0
0
0
9 Inverter~
13 176 119 0 2 22
0 4 20
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
8778 0 0
0
0
9 Inverter~
13 167 84 0 2 22
0 6 21
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
538 0 0
0
0
9 2-In NOR~
219 223 100 0 3 22
0 21 20 19
0
0 0 624 0
6 74LS02
-21 -24 21 -16
3 U1A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 3 2 1 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
6843 0 0
0
0
32
3 1 2 0 0 4240 0 5 8 0 0 3
385 410
435 410
435 407
3 2 3 0 0 8336 0 6 5 0 0 4
282 451
308 451
308 419
333 419
2 1 4 0 0 8336 0 6 1 0 0 3
230 460
97 460
97 71
2 1 5 0 0 4240 0 7 6 0 0 3
200 445
230 445
230 442
1 1 6 0 0 4240 0 2 7 0 0 3
59 70
59 445
164 445
3 1 7 0 0 12432 0 3 5 0 0 4
289 377
308 377
308 401
333 401
0 3 2 0 0 16 0 0 5 0 0 2
380 410
385 410
0 1 6 0 0 16 0 0 3 5 0 4
59 367
58 367
58 368
237 368
0 1 4 0 0 16 0 0 4 3 0 3
97 398
161 398
161 397
2 2 8 0 0 8336 0 4 3 0 0 3
197 397
197 386
237 386
2 1 9 0 0 4224 0 12 9 0 0 3
417 288
436 288
436 285
3 2 10 0 0 8320 0 11 13 0 0 4
283 329
309 329
309 297
334 297
2 0 4 0 0 0 0 11 0 0 3 2
231 338
97 338
2 1 11 0 0 4224 0 10 11 0 0 3
201 323
231 323
231 320
0 1 6 0 0 0 0 0 10 5 0 2
59 323
165 323
3 1 12 0 0 12416 0 15 13 0 0 4
290 255
309 255
309 279
334 279
1 3 13 0 0 4224 0 12 13 0 0 2
381 288
386 288
0 1 6 0 0 0 0 0 15 5 0 3
59 245
59 246
238 246
0 1 4 0 0 0 0 0 14 3 0 3
97 276
162 276
162 275
2 2 14 0 0 8320 0 14 15 0 0 3
198 275
198 264
238 264
0 1 4 0 0 0 0 0 19 3 0 3
97 203
97 202
186 202
0 1 6 0 0 0 0 0 18 5 0 3
59 168
59 167
177 167
2 1 15 0 0 16512 0 16 20 0 0 5
338 166
344 166
344 183
362 183
362 164
3 1 16 0 0 8320 0 17 16 0 0 3
287 183
302 183
302 166
0 1 4 0 0 0 0 0 19 0 0 2
122 202
186 202
2 2 17 0 0 8320 0 19 17 0 0 3
222 202
222 192
235 192
2 1 18 0 0 4224 0 18 17 0 0 4
213 167
225 167
225 174
235 174
1 3 19 0 0 8320 0 21 24 0 0 3
277 92
277 100
262 100
0 1 4 0 0 0 0 0 22 3 0 2
97 119
161 119
0 1 6 0 0 0 0 0 23 5 0 3
59 82
59 84
152 84
2 2 20 0 0 8320 0 22 24 0 0 3
197 119
197 109
210 109
2 1 21 0 0 4224 0 23 24 0 0 4
188 84
200 84
200 91
210 91
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

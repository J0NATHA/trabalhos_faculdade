CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 20 30 100 9
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
100 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 640 259
9961474 0
0
0
0
0
0
0
7
7 Ground~
168 132 154 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
2 +V
167 294 71 0 1 64
0 5
0
0 0 54112 0
3 12V
-11 -13 10 -5
2 V1
-6 -22 8 -14
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
4441 0 0
0
0
11 SPDT Relay~
176 152 98 0 10 64
0 4 6 3 7 2 0 0 0 0
1
0
0 0 864 0
7 12VSPDT
-45 -36 4 -28
4 RLY1
-38 -47 -10 -39
0
0
20 %D %1 %2 %3 %4 %5 %S
0
45 alias:XSPDTRELAY {PULLIN=9.6 RESISTANCE=1000}
4 SIP5
11

0 1 2 3 4 5 1 2 3 4
5 -33686019
88 0 0 0 1 0 0 0
3 RLY
3618 0 0
0
0
11 Signal Gen~
195 40 111 0 24 64
0 7 2 1 86 -7 7 0 0 0
0 0 0 0 0 0 0 1120403456 0 1094713344
0 981668463 981668463 998445679 1008981770
20
0 100 0 12 0 0.001 0.001 0.004 0.01 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
5 0/12V
-17 -28 18 -20
2 V2
-7 -38 7 -30
0
0
40 %D %1 %2 DC 0 PULSE(0 12 0 1m 1m 4m 10m)
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
9 Resistor~
219 209 80 0 4 64
0 4 5 0 1
9 Resistor~
0 0 864 0
2 1k
-10 -13 4 -5
2 R1
-8 -22 6 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
9 Resistor~
219 206 113 0 4 64
0 3 2 0 -1
9 Resistor~
0 0 864 0
3 500
-10 -12 11 -4
2 R2
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7734 0 0
0
0
9 Resistor~
219 215 45 0 4 64
0 6 2 0 -1
9 Resistor~
0 0 864 0
2 1k
-7 -12 7 -4
2 R3
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
9914 0 0
0
0
9
1 3 3 0 0 8320 0 6 3 0 0 4
188 113
174 113
174 87
166 87
1 1 4 0 0 4224 0 3 5 0 0 2
166 80
191 80
2 1 5 0 0 4224 0 5 2 0 0 2
227 80
294 80
2 1 6 0 0 8320 0 3 7 0 0 4
166 73
181 73
181 45
197 45
2 0 2 0 0 8192 0 6 0 0 9 3
224 113
236 113
236 133
4 1 7 0 0 4224 0 3 4 0 0 4
136 93
79 93
79 106
71 106
5 0 2 0 0 0 0 3 0 0 9 3
136 117
119 117
119 133
1 0 2 0 0 0 0 1 0 0 9 2
132 148
132 133
2 2 2 0 0 12416 0 4 7 0 0 6
71 116
89 116
89 133
262 133
262 45
233 45
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.05 0.00025 0.00025
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
2532 8525888 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
0 0 0 0 0 0
16 0
4 0.01 5
1
114 93
0 7 0 0 1	0 6 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

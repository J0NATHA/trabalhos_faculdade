CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 1024 399
7 5.000 V
7 5.000 V
3 GND
1000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 1024 399
9961490 0
0
0
0
0
0
0
11
5 SAVE-
218 309 166 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 B
3 -26 10 -18
5 SAVE1
-11 -36 24 -28
0
0
14 *TRAN -16 32 0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
8953 0 0
0
0
5 SAVE-
218 346 91 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
5 SAVE2
-11 -36 24 -28
0
0
15 *TRAN -54m 15 0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
4441 0 0
0
0
7 Ground~
168 43 154 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
10 Capacitor~
219 43 118 0 2 5
0 3 2
0
0 0 320 270
3 1uF
14 -3 35 5
2 C1
17 -13 31 -5
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
6153 0 0
0
0
2 +V
167 43 81 0 1 3
0 3
0
0 0 53600 0
4 +15V
-12 -16 16 -8
2 V1
-5 -26 9 -18
0
5 DVDD;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
5 4011~
219 301 91 0 3 21
0 4 4 6
0
0 0 96 0
4 4011
-7 -24 21 -16
3 U1B
-4 -34 17 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 2 2 0
1 U
7734 0 0
0
0
5 4011~
219 164 91 0 3 21
0 7 7 4
0
0 0 96 0
4 4011
-7 -24 21 -16
3 U1A
-4 -34 17 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 -1610612720
65 0 0 0 4 1 2 0
1 U
9914 0 0
0
0
4 .IC~
207 239 53 0 1 64
0 4
0
0 0 53568 0
2 0V
-7 -16 7 -8
4 CMD1
-14 -26 14 -18
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 -1610612600
86 0 0 0 1 0 0 0
3 CMD
3747 0 0
0
0
10 Capacitor~
219 355 132 0 2 64
0 6 5
10 Capacitor~
0 0 320 270
5 .01uF
13 -2 48 6
2 C2
21 -15 35 -7
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 -1610612640
67 -1 273 0 1 0 0 0
1 C
3549 0 0
0
0
9 Resistor~
219 227 140 0 2 64
0 5 4
9 Resistor~
0 0 352 90
3 47k
7 -5 28 3
2 R1
10 -15 24 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612600
82 -1 271 0 1 0 0 0
1 R
7931 0 0
0
0
9 Resistor~
219 99 144 0 2 64
0 5 7
9 Resistor~
0 0 352 90
4 470k
8 -5 36 3
2 R2
15 -15 29 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -1610612684
82 -1 271 0 1 0 0 0
1 R
9325 0 0
0
0
11
2 1 2 0 0 4224 0 4 3 0 0 2
43 127
43 148
1 1 3 0 0 4224 0 5 4 0 0 2
43 90
43 109
1 0 4 0 0 4096 0 8 0 0 8 2
239 65
239 91
1 0 5 0 0 4096 0 10 0 0 5 2
227 158
227 166
1 2 5 0 0 8320 0 11 9 0 0 4
99 162
99 166
355 166
355 141
3 1 6 0 0 8320 0 6 9 0 0 3
328 91
355 91
355 123
2 0 4 0 0 4096 0 10 0 0 8 2
227 122
227 91
3 0 4 0 0 4224 0 7 0 0 9 2
191 91
267 91
1 2 4 0 0 0 0 6 6 0 0 4
277 82
267 82
267 100
277 100
2 0 7 0 0 4096 0 7 0 0 11 2
140 100
99 100
2 1 7 0 0 4224 0 11 7 0 0 3
99 126
99 82
140 82
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.005 1e-005 1e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3588 8550976 100 100 0 0
77 66 977 246
0 399 1024 736
977 66
77 66
977 66
977 246
0 0
4.94359e-315 0 5.47077e-315 1.60393e-314 4.94359e-315 4.94359e-315
12409 0
4 0.001 3
1
318 166
0 5 0 0 2	0 5 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
0 66 640 259
9961474 0
0
0
0
0
0
0
5
7 Ground~
168 248 137 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
7 Ground~
168 111 136 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
11 Signal Gen~
195 64 106 0 24 64
0 4 2 1 86 -9 9 0 0 0
0 0 0 0 0 0 0 1268291200 0 1084227584
0 822702175 822702175 850119799 861323157
20
0 2e+007 0 5 0 2e-009 2e-009 2e-008 5e-008 0
0 0 0 0 0 0 0 0 0 0
0
0 0 16976 0
5 -1/1V
-15 -48 20 -40
2 V1
-6 -35 8 -27
0
0
40 %D %1 %2 DC 0 PULSE(0 5 0 2n 2n 20n 50n)
0
0
0
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
13 LossLessLine~
219 173 107 0 4 64
0 4 2 3 2
13 LossLessLine~
0 0 848 0
13 ZO=50 TD=20NS
-46 -20 45 -12
5 LLTR1
-18 -30 17 -22
0
0
17 %D %1 %2 %3 %4 %L
0
0
0
9

0 1 2 3 4 1 2 3 4 -33686019
84 0 0 0 1 0 0 0
4 LLTR
6153 0 0
0
0
9 Resistor~
219 245 103 0 4 64
0 3 2 0 -1
9 Resistor~
0 0 4976 0
2 1k
-7 -12 7 -4
2 R1
-7 -22 7 -14
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
5394 0 0
0
0
6
1 0 2 0 0 4096 0 2 0 0 5 2
111 130
111 111
1 0 2 0 0 4096 0 1 0 0 4 2
248 131
248 111
1 3 3 0 0 4224 0 5 4 0 0 2
227 103
221 103
4 2 2 0 0 4224 0 4 5 0 0 4
221 111
272 111
272 103
263 103
2 2 2 0 0 0 0 3 4 0 0 2
95 111
125 111
1 1 4 0 0 4224 0 4 3 0 0 4
125 103
100 103
100 101
95 101
0
0
16 0 0
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 1e-007 1e-009 1e-009 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
3076 8550464 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
1e-007 0 12 -12 1e-007 1e-007
16 0
4 3e-008 5
1
224 103
0 3 0 0 1	0 3 0 0
0 0 100 100 0 0
98 66 294 126
0 0 0 0
294 66
98 66
294 66
294 126
0 0
1e+007 1 12.16 12.16 1e+007 1e+007
12403 0
0 3e+006 5e+006
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
2000 1 2.36 0 1999 1999
16 0
0 500 1000
0
0 0 100 100 0 0
98 66 296 126
0 0 0 0
296 66
98 66
296 66
296 126
0 0
1e+006 1 -3.55271e-015 -3.55271e-015 999999 999999
12403 0
0 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 644 484
7 5.000 V
7 5.000 V
3 GND
0 66 644 484
135266304 0
0
0
0
0
0
0
17
4 Car~
182 103 316 0 20 64
13 4 6 0 0 0 0 0 0 0
0 0 0 0 4 0 0 0 0 0
400
0
0 0 20528 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 -1610612648
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
9 CA 7-Seg~
184 508 55 0 18 64
10 13 11 12 10 9 8 7 114 3
2 2 2 2 2 2 2 2 1
0
0 0 20512 0
0
0
0
0
0
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 -1610612616
0 0 0 512 1 0 0 0
0
4441 0 0
0
0
9 CA 7-Seg~
184 445 55 0 18 64
10 20 19 18 17 16 15 14 115 3
2 2 2 2 2 2 2 2 1
0
0 0 20512 0
0
0
0
0
0
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 -1610612616
0 0 0 512 1 0 0 0
0
3618 0 0
0
0
9 CA 7-Seg~
184 367 55 0 18 64
10 28 27 26 21 25 24 23 116 3
2 2 2 2 2 2 2 2 1
0
0 0 20512 0
0
0
0
0
0
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 -1610612648
0 0 0 512 1 0 0 0
0
6153 0 0
0
0
9 CA 7-Seg~
184 304 55 0 18 64
10 34 33 32 22 31 30 29 117 3
2 2 2 2 2 2 2 2 1
0
0 0 20512 0
0
0
0
0
0
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 -1610612616
0 0 0 512 1 0 0 0
0
5394 0 0
0
0
4 Car~
182 103 278 0 20 64
12 4 35 0 0 0 0 0 0 0
0 0 0 0 3 0 0 0 0 0
400
0
0 0 20528 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 -1610612616
0 0 0 0 1 0 0 0
0
7734 0 0
0
0
4 Car~
182 104 240 0 20 64
10 4 36 0 0 0 0 0 0 0
0 0 0 0 4 0 0 0 0 0
400
0
0 0 20528 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 -1610612616
0 0 0 0 1 0 0 0
0
9914 0 0
0
0
7 Pulser~
4 63 153 0 10 64
0 118 119 5 120 0 0 5 5 2
7
0
0 0 20528 0
0
0
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 -1610612616
0 0 0 512 1 0 0 0
0
3747 0 0
0
0
7 Ground~
168 13 265 0 1 64
0 2
0
0 0 53360 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -1610612487
0 0 0 0 1 0 0 0
0
3549 0 0
0
0
14 NO PushButton~
191 48 85 0 2 64
0 3 4
0
0 0 20592 0
0
0
0
0
0
0
0
0
5

0 1 2 1 2 -1610612616
0 0 0 0 1 0 0 0
1 S
7931 0 0
0
0
2 +V
167 82 24 0 1 64
0 3
0
0 0 53488 0
3 10V
-10 -22 11 -14
0
0
4 VCC;
10 %D %1 0 %V
0
0
0
3

0 1 1 -1610612616
86 0 0 0 1 0 0 0
1 V
9325 0 0
0
0
9 CA 7-Seg~
184 229 54 0 18 64
10 46 47 48 49 45 44 43 121 3
2 2 2 2 2 2 2 2 1
0
0 0 20512 0
0
0
0
0
0
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 -1610612616
0 0 0 512 1 0 0 0
0
8903 0 0
0
0
9 CA 7-Seg~
184 166 54 0 18 64
10 37 38 39 50 42 41 40 122 3
2 2 2 2 2 2 2 2 1
0
0 0 20512 0
0
0
0
0
0
0
0
0
19

0 1 2 3 4 5 6 7 8 9
1 2 3 4 5 6 7 8 9 -1610612632
0 0 0 512 1 0 0 0
0
3834 0 0
0
0
6 Timer~
94 199 148 0 17 64
0 44 45 49 48 47 46 40 41 42
50 39 38 37 43 5 4 36
6 Timer~
1 0 4528 90
7 Red Car
-33 -3 16 5
0
0
0
0
0
0
0
35

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 -1610612712
0 0 0 0 1 0 0 0
1 U
3363 0 0
0
0
6 Timer~
94 337 148 0 17 64
0 24 25 21 26 27 28 29 30 31
22 32 33 34 23 5 4 35
6 Timer~
2 0 4528 90
9 Green Car
-37 -3 26 5
0
0
0
0
0
0
0
35

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 -1610612632
0 0 0 0 1 0 0 0
1 U
7668 0 0
0
0
6 Timer~
94 478 148 0 17 64
0 8 9 10 12 11 13 14 15 16
17 18 19 20 7 5 4 6
6 Timer~
3 0 4528 90
8 Blue Car
-35 -2 21 6
0
0
0
0
0
0
0
35

0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0 0 0 0 0 -1610612632
0 0 0 0 1 0 0 0
1 U
4718 0 0
0
0
9 Resistor~
219 13 229 0 3 64
0 2 4 -1
9 Resistor~
0 0 4208 90
2 1k
-7 -28 7 -20
0
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 -1610612495
82 0 0 0 1 0 0 0
1 R
3874 0 0
0
0
63
1 1 2 0 0 4224 0 9 17 0 0 2
13 259
13 247
1 0 4 0 0 4096 0 7 0 0 4 2
64 235
29 235
1 0 4 0 0 0 0 6 0 0 4 2
63 273
29 273
0 1 4 0 0 4096 0 0 1 44 0 3
29 197
29 311
63 311
15 0 5 0 0 4224 0 16 0 0 42 2
427 185
286 185
2 17 6 0 0 12416 0 1 16 0 0 5
63 320
57 320
57 226
445 226
445 179
0 16 4 0 0 4096 0 0 16 41 0 3
295 197
436 197
436 179
7 14 7 0 0 12416 0 2 16 0 0 4
523 91
523 98
529 98
529 115
1 6 8 0 0 4224 0 16 2 0 0 4
521 115
521 103
517 103
517 91
5 2 9 0 0 4224 0 2 16 0 0 4
511 91
511 108
513 108
513 115
3 4 10 0 0 4224 0 16 2 0 0 2
505 115
505 91
2 5 11 0 0 4224 0 2 16 0 0 4
493 91
493 103
489 103
489 115
3 4 12 0 0 4224 0 2 16 0 0 4
499 91
499 108
497 108
497 115
1 6 13 0 0 12416 0 2 16 0 0 4
487 91
487 98
480 98
480 115
9 0 3 0 0 4096 0 3 0 0 16 2
445 19
445 9
0 9 3 0 0 4224 0 0 2 39 0 3
367 9
508 9
508 19
7 7 14 0 0 12416 0 3 16 0 0 4
460 91
460 98
467 98
467 115
6 8 15 0 0 4224 0 3 16 0 0 4
454 91
454 103
459 103
459 115
5 9 16 0 0 4224 0 3 16 0 0 4
448 91
448 108
450 108
450 115
10 4 17 0 0 4224 0 16 3 0 0 2
442 115
442 91
3 11 18 0 0 4224 0 3 16 0 0 4
436 91
436 108
434 108
434 115
2 12 19 0 0 4224 0 3 16 0 0 4
430 91
430 103
426 103
426 115
1 13 20 0 0 12416 0 3 16 0 0 4
424 91
424 98
418 98
418 115
3 4 21 0 0 4224 0 15 4 0 0 2
364 115
364 91
10 4 22 0 0 4224 0 15 5 0 0 2
301 115
301 91
7 14 23 0 0 12416 0 4 15 0 0 4
382 91
382 98
388 98
388 115
6 1 24 0 0 4224 0 4 15 0 0 4
376 91
376 103
380 103
380 115
5 2 25 0 0 4224 0 4 15 0 0 4
370 91
370 108
372 108
372 115
3 4 26 0 0 4224 0 4 15 0 0 4
358 91
358 108
356 108
356 115
5 2 27 0 0 4224 0 15 4 0 0 4
348 115
348 103
352 103
352 91
1 6 28 0 0 12416 0 4 15 0 0 4
346 91
346 98
339 98
339 115
7 7 29 0 0 4224 0 5 15 0 0 4
319 91
319 103
326 103
326 115
6 8 30 0 0 4224 0 5 15 0 0 4
313 91
313 103
318 103
318 115
5 9 31 0 0 4224 0 5 15 0 0 4
307 91
307 108
309 108
309 115
3 11 32 0 0 4224 0 5 15 0 0 4
295 91
295 108
293 108
293 115
2 12 33 0 0 4224 0 5 15 0 0 4
289 91
289 103
285 103
285 115
1 13 34 0 0 12416 0 5 15 0 0 4
283 91
283 98
277 98
277 115
9 0 3 0 0 0 0 5 0 0 39 2
304 19
304 9
0 9 3 0 0 0 0 0 4 47 0 3
229 9
367 9
367 19
2 17 35 0 0 12416 0 6 15 0 0 5
63 282
48 282
48 216
304 216
304 179
0 16 4 0 0 0 0 0 15 44 0 3
157 197
295 197
295 179
15 15 5 0 0 0 0 14 15 0 0 2
148 185
286 185
2 17 36 0 0 12416 0 7 14 0 0 5
64 244
38 244
38 207
166 207
166 179
16 0 4 0 0 8320 0 14 0 0 49 3
157 179
157 197
13 197
3 15 5 0 0 0 0 8 14 0 0 4
87 144
112 144
112 185
148 185
9 0 3 0 0 0 0 13 0 0 47 2
166 18
166 9
9 0 3 0 0 0 0 12 0 0 48 5
229 18
229 9
127 9
127 46
82 46
1 1 3 0 0 0 0 10 11 0 0 3
65 93
82 93
82 33
2 2 4 0 0 0 0 10 17 0 0 3
31 93
13 93
13 211
1 13 37 0 0 12416 0 13 14 0 0 4
145 90
145 98
139 98
139 115
2 12 38 0 0 4224 0 13 14 0 0 4
151 90
151 103
147 103
147 115
3 11 39 0 0 4224 0 13 14 0 0 4
157 90
157 108
155 108
155 115
7 7 40 0 0 12416 0 13 14 0 0 4
181 90
181 98
188 98
188 115
6 8 41 0 0 4224 0 13 14 0 0 4
175 90
175 103
180 103
180 115
5 9 42 0 0 4224 0 13 14 0 0 4
169 90
169 108
171 108
171 115
7 14 43 0 0 12416 0 12 14 0 0 4
244 90
244 98
250 98
250 115
6 1 44 0 0 4224 0 12 14 0 0 4
238 90
238 103
242 103
242 115
5 2 45 0 0 4224 0 12 14 0 0 4
232 90
232 108
234 108
234 115
1 6 46 0 0 12416 0 12 14 0 0 4
208 90
208 98
201 98
201 115
2 5 47 0 0 4224 0 12 14 0 0 4
214 90
214 103
210 103
210 115
3 4 48 0 0 4224 0 12 14 0 0 4
220 90
220 108
218 108
218 115
3 4 49 0 0 4224 0 14 12 0 0 2
226 115
226 90
4 10 50 0 0 4224 0 13 14 0 0 2
163 90
163 115
1
16 8 0 0 0 0 0 0 0 0 0 0 54
6 System
0 0 0 5
29 98 73 120
33 102 63 118
5 Start
0
0 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 71 1536 816
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
80 C:\Users\jonat\AppData\Local\Temp\Rar$EXa10028.42639\CIRCUIT MAKER_CM60S\BOM.DAT
0 7
0 71 1536 816
143654930 0
0
6 Title:
5 Name:
0
0
0
35
13 Logic Switch~
5 99 37 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 74 37 0 1 11
0 5
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
9 Inverter~
13 415 479 0 2 22
0 3 2
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U7A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 7 0
1 U
3618 0 0
0
0
9 Inverter~
13 214 456 0 2 22
0 13 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 5 0
1 U
6153 0 0
0
0
10 2-In NAND~
219 172 456 0 3 22
0 11 4 13
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U6A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
5394 0 0
0
0
10 2-In NAND~
219 169 503 0 3 22
0 5 10 12
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U4D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 4 0
1 U
7734 0 0
0
0
9 Inverter~
13 211 503 0 2 22
0 12 7
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 5 0
1 U
9914 0 0
0
0
9 Inverter~
13 121 447 0 2 22
0 5 11
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 5 0
1 U
3747 0 0
0
0
9 Inverter~
13 126 529 0 2 22
0 4 10
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 5 0
1 U
3549 0 0
0
0
9 Inverter~
13 315 513 0 2 22
0 7 8
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 5 0
1 U
7931 0 0
0
0
9 Inverter~
13 301 457 0 2 22
0 6 9
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U5A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 5 0
1 U
9325 0 0
0
0
10 2-In NAND~
219 370 477 0 3 22
0 9 8 3
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U4C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 4 0
1 U
8903 0 0
0
0
14 Logic Display~
6 451 457 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3834 0 0
0
0
14 Logic Display~
6 423 325 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3363 0 0
0
0
10 2-In NAND~
219 371 345 0 3 22
0 17 16 18
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U4B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 4 0
1 U
7668 0 0
0
0
9 Inverter~
13 302 325 0 2 22
0 14 17
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 3 0
1 U
4718 0 0
0
0
9 Inverter~
13 316 381 0 2 22
0 15 16
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 3 0
1 U
3874 0 0
0
0
9 Inverter~
13 127 397 0 2 22
0 4 19
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 3 0
1 U
6671 0 0
0
0
9 Inverter~
13 122 315 0 2 22
0 5 20
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 3 0
1 U
3789 0 0
0
0
9 Inverter~
13 212 371 0 2 22
0 21 15
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 3 0
1 U
4871 0 0
0
0
10 2-In NAND~
219 170 371 0 3 22
0 5 19 21
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U4A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3750 0 0
0
0
10 2-In NAND~
219 173 324 0 3 22
0 20 4 22
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1D
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 4 1 0
1 U
8778 0 0
0
0
9 Inverter~
13 215 324 0 2 22
0 22 14
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U3A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 3 0
1 U
538 0 0
0
0
9 Inverter~
13 261 242 0 2 22
0 24 23
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2B
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 2 0
1 U
6843 0 0
0
0
14 Logic Display~
6 298 223 0 1 2
10 23
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3136 0 0
0
0
10 2-In NAND~
219 211 242 0 3 22
0 26 25 24
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1C
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 10 9 8 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 3 1 0
1 U
5950 0 0
0
0
9 Inverter~
13 144 231 0 2 22
0 5 26
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2F
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 6 2 0
1 U
5670 0 0
0
0
9 Inverter~
13 149 277 0 2 22
0 4 25
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2E
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 5 2 0
1 U
6828 0 0
0
0
9 Inverter~
13 158 187 0 2 22
0 4 27
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2D
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 4 2 0
1 U
6735 0 0
0
0
9 Inverter~
13 144 131 0 2 22
0 5 28
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2C
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 2 0
1 U
8365 0 0
0
0
10 2-In NAND~
219 213 151 0 3 22
0 28 27 29
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
4132 0 0
0
0
14 Logic Display~
6 265 131 0 1 2
10 29
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4551 0 0
0
0
14 Logic Display~
6 251 55 0 1 2
10 30
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3635 0 0
0
0
9 Inverter~
13 217 74 0 2 22
0 31 30
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 U2A
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 1 2 0
1 U
3973 0 0
0
0
10 2-In NAND~
219 175 74 0 3 22
0 5 4 31
0
0 0 624 0
6 74LS00
-14 -24 28 -16
3 U1A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
3851 0 0
0
0
46
1 2 2 0 0 8320 0 13 3 0 0 4
451 475
451 478
436 478
436 479
1 3 3 0 0 4224 0 3 12 0 0 4
400 479
394 479
394 477
397 477
1 0 4 0 0 4096 0 9 0 0 45 2
111 529
99 529
1 0 5 0 0 4096 0 8 0 0 46 2
106 447
74 447
2 0 6 0 0 4096 0 4 0 0 7 2
235 456
235 457
1 2 7 0 0 4224 0 10 7 0 0 4
300 513
258 513
258 503
232 503
1 0 6 0 0 4224 0 11 0 0 0 2
286 457
231 457
2 2 8 0 0 8320 0 10 12 0 0 5
336 513
339 513
339 495
346 495
346 486
2 1 9 0 0 4224 0 11 12 0 0 3
322 457
346 457
346 468
2 2 10 0 0 8320 0 9 6 0 0 4
147 529
144 529
144 512
145 512
2 1 11 0 0 4224 0 8 5 0 0 2
142 447
148 447
1 0 5 0 0 4096 0 6 0 0 46 2
145 494
74 494
1 3 12 0 0 0 0 7 6 0 0 2
196 503
196 503
2 0 4 0 0 4096 0 5 0 0 45 2
148 465
99 465
1 3 13 0 0 0 0 4 5 0 0 2
199 456
199 456
2 0 14 0 0 4096 0 23 0 0 18 2
236 324
236 325
1 2 15 0 0 4224 0 17 20 0 0 4
301 381
259 381
259 371
233 371
1 0 14 0 0 4224 0 16 0 0 0 2
287 325
232 325
2 2 16 0 0 8320 0 17 15 0 0 5
337 381
340 381
340 363
347 363
347 354
2 1 17 0 0 4224 0 16 15 0 0 3
323 325
347 325
347 336
1 3 18 0 0 8320 0 14 15 0 0 5
423 343
423 344
399 344
399 345
398 345
2 2 19 0 0 8320 0 18 21 0 0 4
148 397
145 397
145 380
146 380
2 1 20 0 0 4224 0 19 22 0 0 2
143 315
149 315
0 1 4 0 0 0 0 0 18 45 0 4
99 380
103 380
103 397
112 397
1 0 5 0 0 4096 0 21 0 0 46 2
146 362
74 362
1 3 21 0 0 0 0 20 21 0 0 2
197 371
197 371
2 0 4 0 0 4096 0 22 0 0 45 2
149 333
99 333
0 1 5 0 0 0 0 0 19 46 0 2
74 315
107 315
1 3 22 0 0 0 0 23 22 0 0 2
200 324
200 324
2 1 23 0 0 4224 0 24 25 0 0 3
282 242
298 242
298 241
1 0 4 0 0 0 0 28 0 0 45 2
134 277
99 277
1 0 4 0 0 0 0 29 0 0 45 2
143 187
99 187
2 0 4 0 0 4096 0 35 0 0 45 2
151 83
99 83
3 1 24 0 0 4224 0 26 24 0 0 2
238 242
246 242
1 0 5 0 0 0 0 27 0 0 46 2
129 231
74 231
2 2 25 0 0 8320 0 28 26 0 0 3
170 277
187 277
187 251
2 1 26 0 0 8320 0 27 26 0 0 4
165 231
165 234
187 234
187 233
1 0 5 0 0 0 0 30 0 0 46 2
129 131
74 131
2 2 27 0 0 8320 0 29 31 0 0 5
179 187
182 187
182 169
189 169
189 160
2 1 28 0 0 4224 0 30 31 0 0 3
165 131
189 131
189 142
1 3 29 0 0 8320 0 32 31 0 0 5
265 149
265 150
241 150
241 151
240 151
1 2 30 0 0 8320 0 33 34 0 0 3
251 73
251 74
238 74
1 0 5 0 0 4096 0 35 0 0 46 2
151 65
74 65
1 3 31 0 0 0 0 34 35 0 0 2
202 74
202 74
1 0 4 0 0 4224 0 1 0 0 0 2
99 49
99 602
1 0 5 0 0 4224 0 2 0 0 0 2
74 49
74 603
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

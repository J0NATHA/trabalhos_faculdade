CircuitMaker Text
4
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 1e+012
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 0
0 66 240 382
0 66 240 382
9961474 0
0
0
0
0
0
0
9
5 SAVE-
218 105 163 0 11 
0 0 0 0 0 0 0 0 0 0 
1 0 0
0 0 -8000 0
1 B
3 -26 10 -18
0
0
0
12 *TRAN 0 5.76
0
1

0 0 
0 0 0 0 0 0 0 0
0
8953 0 0 0
5 SAVE-
218 67 128 0 11 
0 0 0 0 0 0 0 0 0 0 
1 0 0
0 0 -8000 0
1 A
3 -26 10 -18
0
0
0
12 *TRAN 0 11.7
0
1

0 0 
0 0 0 0 0 0 0 0
0
4441 0 0 0
2 +V
167 75 32 0 2 
0 6 0 0
0 0 -11936 0
3 20V
-10 -14 11 -6
2 V1
-7 -24 7 -16
0
0
13 %D %1 0 DC %V
0
2

0 1 0 
86 0 0 0 0 0 0 0
1 V
3618 0 0 0
7 Ground~
168 75 237 0 2 
0 2 0 0
0 0 -12192 0
0
0
0
4 GND;
0
0
2

0 1 0 
0 0 0 0 0 0 0 0
0
6153 0 0 0
6 N-UJT~
94 97 136 0 4 
0 5 3 4 0 6 N-UJT~
1 0 320 0
6 2N2646
6 -3 48 5
2 Q1
20 -13 34 -5
0
0
14 %D %1 %2 %3 %S
0
4

0 1 2 3 0 
88 0 0 0 0 0 0 0
1 Q
5394 0 0 0
10 Capacitor~
94 49 173 0 3 
0 2 5 0 10 Capacitor~
2 0 320 90
4 .1uF
-39 -3 -11 5
2 C1
-32 -13 -18 -5
6 CAP0.2
-22 -38 20 -30
0
11 %D %1 %2 %V
0
3

0 1 2 0 
67 0 0 0 0 0 0 0
1 C
7734 0 0 0
9 Resistor~
94 105 186 0 4 
0 2 3 -1 0 9 Resistor~
3 0 4448 90
2 47
11 -2 25 6
2 R1
11 -12 25 -4
0
0
11 %D %1 %2 %V
0
3

0 1 2 0 
82 0 0 0 0 0 0 0
1 R
9914 0 0 0
9 Resistor~
94 105 88 0 5 
0 4 6 0 1 0 9 Resistor~
4 0 4448 90
3 330
7 2 28 10
2 R2
10 -8 24 0
0
0
11 %D %1 %2 %V
0
3

0 1 2 0 
82 0 0 0 0 0 0 0
1 R
3747 0 0 0
9 Resistor~
94 49 90 0 5 
0 5 6 0 1 0 9 Resistor~
5 0 4448 90
3 50k
-26 -1 -5 7
2 R3
-18 -11 -4 -3
0
0
11 %D %1 %2 %V
0
3

0 1 2 0 
82 0 0 0 0 0 0 0
1 R
3549 0 0 0
8
2 2 3 0 0 4224 0 5 7 0 0 2
105 154
105 168
3 1 4 0 0 4224 0 5 8 0 0 2
105 118
105 106
1 0 5 0 0 4096 0 5 0 0 8 2
83 128
49 128
1 0 6 0 0 4096 0 3 0 0 7 2
75 41
75 58
1 0 2 0 0 4096 0 4 0 0 6 2
75 231
75 215
1 1 2 0 0 8320 0 7 6 0 0 4
105 204
105 215
49 215
49 182
2 2 6 0 0 8320 0 8 9 0 0 4
105 70
105 58
49 58
49 72
1 2 5 0 0 4224 0 9 6 0 0 2
49 108
49 164
0
0
16 2 0
0
0
0
0 0 0
0
0 0 0
0 0 1 2
0 0.015 0.0001 0.0001 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

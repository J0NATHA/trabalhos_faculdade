CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 3
0 66 640 259
7 5.000 V
7 5.000 V
3 GND
0 66 640 259
144179216 0
0
0
0
0
0
0
8
5 SAVE-
218 138 19 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
16 *DC 872n 8.63m 0
0
0
0
11

0 0 0 0 0 0 0 0 0 0
0 0
0 0 0 0 1 0 0 0
4 SAVE
8953 0 0
0
0
9 I Source~
198 67 113 0 2 5
0 4 2
0
0 0 16992 0
5 100mA
12 -2 47 6
3 Ibb
19 -12 40 -4
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
73 0 0 0 0 0 0 0
2 Is
4441 0 0
0
0
9 V Source~
197 250 61 0 2 5
0 5 2
0
0 0 16992 0
3 10V
12 -2 33 6
3 Vce
12 -12 33 -4
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
3618 0 0
0
0
9 V Source~
197 138 37 0 2 5
0 5 3
0
0 0 16736 0
2 0V
15 -2 29 6
3 Vs1
12 -12 33 -4
0
0
11 %D %1 %2 %V
0
0
0
5

0 1 2 1 2 0
86 0 0 0 0 0 0 0
2 Vs
6153 0 0
0
0
7 Ground~
168 250 118 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
5394 0 0
0
0
7 Ground~
168 67 149 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7734 0 0
0
0
7 Ground~
168 138 128 0 1 3
0 2
0
0 0 53344 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
9914 0 0
0
0
12 PNP Trans:C~
219 133 86 0 3 7
0 2 4 3
12 NPN Trans:C~
0 0 320 692
6 2N3906
20 -4 62 4
2 Q1
33 -14 47 -6
0
0
14 %D %1 %2 %3 %M
0
0
6 TO-92B
7

0 1 2 3 1 2 3 -33686019
113 -1 261 0 1 1 0 0
1 Q
3747 0 0
0
0
6
1 1 2 0 0 4096 0 8 7 0 0 2
138 104
138 122
2 3 3 0 0 4224 0 4 8 0 0 2
138 58
138 68
2 1 4 0 0 4224 0 8 2 0 0 3
115 86
67 86
67 92
2 1 2 0 0 0 0 2 6 0 0 2
67 134
67 143
1 1 5 0 0 8320 0 3 4 0 0 4
250 40
250 8
138 8
138 16
2 1 2 0 0 4224 0 3 5 0 0 2
250 82
250 112
0
0
4 0 0
0
0
3 Vce
0 4 0.02
3 Ibb
1e-005 8e-005 1e-005
3 0 1 4
0 2e-006 1e-008 1e-008 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
2052 2259008 100 100 0 0
77 66 617 126
0 259 640 452
617 66
77 66
617 66
617 126
0 0
5.34602e-315 0 4.99564e-315 0 5.34602e-315 4.99564e-315
0 0
4 1 3
1
138 19
0 5 0 0 1	4 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 66 1024 399
8  5.000 V
8  5.000 V
3 GND
500 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 1024 399
9961490 0
0
0
0
0
0
0
9
5 SAVE-
218 236 105 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
5 SAVE1
-11 -36 24 -28
0
0
12 *TRAN 0 12 0
0
0
0
3

0 0 0 0
0 0 0 0 1 0 0 0
4 SAVE
8953 0 0
0
0
4 .IC~
207 186 76 0 1 3
0 4
0
0 0 53568 0
2 0V
-7 -16 7 -8
4 CMD1
-14 -26 14 -18
0
0
12 .IC V(%1)=%V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
3 CMD
4441 0 0
0
0
7 Ground~
168 268 185 0 1 3
0 2
0
0 0 53344 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3618 0 0
0
0
7 Ground~
168 186 224 0 1 3
0 2
0
0 0 53344 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6153 0 0
0
0
2 +V
167 88 56 0 1 3
0 3
0
0 0 54624 0
4 +12V
-13 -14 15 -6
2 V1
-7 -32 7 -24
3 VDD
-9 -26 12 -18
5 DVDD;
13 %D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 0 0
1 V
5394 0 0
0
0
10 Capacitor~
219 186 196 0 2 5
0 5 2
0
0 0 320 270
3 1uF
11 -5 32 3
2 C1
14 -15 28 -7
0
0
11 %D %1 %2 %V
0
0
6 RAD0.2
5

0 1 2 1 2 0
67 0 0 0 1 0 0 0
1 C
7734 0 0
0
0
5 4093~
219 119 105 0 3 21
0 3 5 4
0
0 0 352 0
4 4093
2 -26 30 -18
3 U1A
-4 -34 17 -26
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
16

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0
65 0 0 0 4 1 1 0
1 U
9914 0 0
0
0
9 Resistor~
219 268 138 0 4 5
0 4 2 0 -1
0
0 0 352 270
3 27k
5 -5 26 3
2 R1
8 -15 22 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 186 141 0 2 5
0 4 5
0
0 0 352 270
2 1k
8 -5 22 3
2 R2
8 -15 22 -7
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 0
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
8
1 0 4 0 0 4096 0 2 0 0 7 2
186 88
186 105
1 2 2 0 0 4096 0 4 6 0 0 2
186 218
186 205
1 2 2 0 0 4224 0 3 8 0 0 2
268 179
268 156
0 2 5 0 0 4224 0 0 7 5 0 4
186 172
87 172
87 114
95 114
2 1 5 0 0 0 0 9 6 0 0 2
186 159
186 187
1 0 4 0 0 4096 0 9 0 0 7 2
186 123
186 105
3 1 4 0 0 4224 0 7 8 0 0 3
146 105
268 105
268 120
1 1 3 0 0 4224 0 5 7 0 0 3
88 65
88 96
95 96
0
0
16 0 1
0
0
0
0 0 0
0
0 0 0
3 0 1 4
0 0.01 1e-005 1e-005
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3084 8550976 100 100 0 0
77 66 977 246
0 399 1024 736
977 66
77 66
977 66
977 246
0 0
4.98503e-315 0 5.4086e-315 0 4.98503e-315 4.98503e-315
12409 0
4 0.003 2
1
257 105
0 4 0 0 1	0 7 0 0
3688 8550464 100 100 0 0
77 66 977 276
0 403 1024 740
977 66
77 66
977 66
977 276
0 0
0 0 0 0 0 0
16 0
4 1e-006 2
1
343 149
0 3 0 0 1	0 9 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

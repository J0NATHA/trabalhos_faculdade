CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 10 100 9
0 66 320 259
7 5.000 V
7 5.000 V
3 GND
10000 10
24 100 1 1 0
20 Package,Description,
18 C:\CM50_32\BOM.DAT
0 7
0 66 320 259
12058632 1
0
0
0
0
0
0
10
5 SAVE-
218 199 70 0 10 11
0 0 0 0 0 0 0 0 0 0
1
0
0 0 57536 0
1 A
3 -26 10 -18
0
0
0
10 *TRAN -1 1
0
0
0
3

0 0 0 -33686019
0 0 0 0 1 0 0 0
0
8953 0 0
0
0
7 Ground~
168 198 158 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
4441 0 0
0
0
2 +V
167 153 135 0 1 64
0 4
0
0 0 54112 180
4 -12V
-14 0 14 8
3 Vee
-9 10 12 18
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
3618 0 0
0
0
2 +V
167 153 59 0 1 64
0 3
0
0 0 54112 0
4 +12v
-13 -13 15 -5
3 Vcc
-9 -23 12 -15
0
0
13 %D %1 0 DC %V
0
0
0
3

0 1 1 -33686019
86 0 0 0 1 0 0 0
1 V
6153 0 0
0
0
7 Ground~
168 101 131 0 1 64
0 2
0
0 0 53344 0
0
0
0
4 GND;
0
0
0
0
3

0 1 1 -33686019
0 0 0 0 1 0 0 0
0
5394 0 0
0
0
11 Signal Gen~
195 41 93 0 19 64
0 7 2 2 86 -8 8 0 0 0
0 0 0 0 0 0 -1110651699 1176256512 0 1036831949
20
-0.1 10000 0 0.1 0 0 0 0 0 0
0 0 0 0 0 0 0 0 0 0
0
0 0 832 0
11 -100m/100mV
-38 23 39 31
3 Vin
-11 -31 10 -23
0
0
44 %D %1 %2 DC 0 SIN(0 100m 10k 0 0) AC -100m 0
0
0
4 SIP2
5

0 1 2 1 2 -33686019
86 0 0 0 1 0 0 0
1 V
7734 0 0
0
0
8 Op-Amp5~
219 153 94 0 5 64
0 2 5 3 4 6
8 Op-Amp5~
0 0 832 0
5 UA741
7 -13 42 -5
2 U1
15 -23 29 -15
0
0
20 %D %1 %2 %3 %4 %5 %S
0
0
4 DIP8
11

0 3 2 7 4 6 3 2 7 4
6 -33686019
88 0 0 0 1 0 0 0
1 U
9914 0 0
0
0
9 Resistor~
219 101 88 0 2 64
0 7 5
9 Resistor~
0 0 4960 0
3 10k
-10 -12 11 -4
2 RI
-6 -23 8 -15
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3747 0 0
0
0
9 Resistor~
219 164 25 0 2 64
0 5 6
9 Resistor~
0 0 4960 0
6 100.0k
-20 -12 22 -4
2 RF
-6 -22 8 -14
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
3549 0 0
0
0
9 Resistor~
219 198 122 0 3 64
0 2 6 -1
9 Resistor~
0 0 4960 90
3 25k
5 1 26 9
2 RL
7 -9 21 -1
0
0
11 %D %1 %2 %V
0
0
8 AXIAL0.4
5

0 1 2 1 2 -33686019
82 0 0 0 1 0 0 0
1 R
7931 0 0
0
0
10
1 0 2 0 0 4096 0 5 0 0 2 2
101 125
101 100
1 2 2 0 0 4224 0 7 6 0 0 4
135 100
83 100
83 98
72 98
1 1 2 0 0 0 0 10 2 0 0 2
198 140
198 152
3 1 3 0 0 4224 0 7 4 0 0 2
153 81
153 68
4 1 4 0 0 4224 0 7 3 0 0 2
153 107
153 120
1 0 5 0 0 8320 0 9 0 0 7 3
146 25
127 25
127 88
2 2 5 0 0 0 0 8 7 0 0 2
119 88
135 88
2 0 6 0 0 8320 0 9 0 0 9 3
182 25
198 25
198 94
5 2 6 0 0 0 0 7 10 0 0 3
171 94
198 94
198 104
1 1 7 0 0 4224 0 6 8 0 0 2
72 88
83 88
0
0
29 0 1
0
0
3 Vin
-0.7 -1.5 -0.02
0
0 0 0
100 0 1 1e+006
0 0.0005 2.5e-006 2.5e-006
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
3236 1210432 100 100 0 0
77 66 617 126
0 66 140 136
617 66
77 66
617 66
617 126
0 0
4.80864e-315 0 5.27183e-315 1.58818e-314 4.80864e-315 5.31328e-315
16 0
4 1 5
1
153 76
0 3 0 0 1	0 4 0 0
756 8550464 100 100 0 0
77 66 287 126
0 259 320 452
286 66
77 66
287 66
287 126
0 0
4.80864e-315 0 5.27183e-315 1.58818e-314 4.80864e-315 4.80864e-315
16 0
4 0.0001 5
2
78 88
0 7 0 0 1	0 10 0 0
198 60
0 6 0 0 2	0 8 0 0
3552 2259008 100 100 0 0
77 66 287 126
320 66 640 259
287 66
77 66
287 66
287 126
0 0
1.58487e-314 1.58934e-314 5.39928e-315 5.37337e-315 5.24531e-315 5.24531e-315
0 0
4 0.3 5
1
198 62
0 6 0 0 2	0 8 0 0
3600 4421696 100 100 0 0
98 66 296 126
320 259 640 452
296 66
98 66
296 66
296 66
0 0
6.08861e-315 5.26354e-315 1.38842e-314 0 6.08861e-315 6.08861e-315
12403 0
4 300000 500000
1
198 67
0 6 0 0 2	0 8 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

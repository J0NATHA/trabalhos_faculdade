CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
20 81 1480 777
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
80 C:\Users\jonat\AppData\Local\Temp\Rar$EXa47972.16692\CIRCUIT MAKER_CM60S\BOM.DAT
0 7
20 81 1480 777
143654930 0
0
6 Title:
5 Name:
0
0
0
11
13 Logic Switch~
5 183 62 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 154 61 0 10 11
0 9 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 120 61 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -22 8 -14
1 A
-3 -32 4 -24
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
3618 0 0
0
0
9 Inverter~
13 285 155 0 2 22
0 4 3
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 NOC
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 3 4 0
1 U
6153 0 0
0
0
9 Inverter~
13 294 84 0 2 22
0 7 6
0
0 0 624 0
6 74LS04
-21 -19 21 -11
3 NOB
-11 -20 10 -12
0
15 DVCC=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 0 0
65 0 0 0 6 2 4 0
1 U
5394 0 0
0
0
9 2-In XOR~
219 220 252 0 3 22
0 9 8 5
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 XOB
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
7734 0 0
0
0
9 2-In AND~
219 333 203 0 3 22
0 4 5 2
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 ANB
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 2 0
1 U
9914 0 0
0
0
14 Logic Display~
6 465 158 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3747 0 0
0
0
8 2-In OR~
219 394 160 0 3 22
0 11 2 10
0
0 0 624 0
6 74LS32
-21 -24 21 -16
2 OR
0 -25 14 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 3 0
1 U
3549 0 0
0
0
9 2-In AND~
219 336 118 0 3 22
0 6 3 11
0
0 0 624 0
6 74LS08
-21 -24 21 -16
3 AND
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7931 0 0
0
0
9 2-In XOR~
219 247 115 0 3 22
0 9 8 7
0
0 0 624 0
6 74LS86
-21 -24 21 -16
3 XOR
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 1 0
1 U
9325 0 0
0
0
16
3 2 2 0 0 8320 0 7 9 0 0 4
354 203
373 203
373 169
381 169
2 2 3 0 0 8336 0 4 10 0 0 4
306 155
311 155
311 127
312 127
0 1 4 0 0 4096 0 0 4 16 0 3
120 148
270 148
270 155
0 1 4 0 0 4096 0 0 7 16 0 2
120 194
309 194
2 3 5 0 0 8320 0 7 6 0 0 3
309 212
309 252
253 252
1 2 6 0 0 8320 0 10 5 0 0 4
312 109
313 109
313 84
315 84
1 3 7 0 0 4224 0 5 11 0 0 3
279 84
279 115
280 115
0 2 8 0 0 4096 0 0 6 15 0 3
183 222
183 261
204 261
0 1 9 0 0 8192 0 0 6 14 0 3
154 202
154 243
204 243
3 1 10 0 0 8320 0 9 8 0 0 5
427 160
442 160
442 188
465 188
465 176
3 1 11 0 0 8320 0 10 9 0 0 4
357 118
369 118
369 151
381 151
0 2 8 0 0 4096 0 0 11 15 0 2
183 124
231 124
0 1 9 0 0 8192 0 0 11 14 0 3
154 105
154 106
231 106
1 0 9 0 0 4224 0 2 0 0 0 2
154 73
154 420
1 0 8 0 0 4224 0 1 0 0 0 2
183 74
183 422
1 0 4 0 0 4224 0 3 0 0 0 2
120 73
120 419
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

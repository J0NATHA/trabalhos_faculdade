CircuitMaker Text
5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 19 14 16 20 20 20 20 10 13 
20 18 11 
0 0 3 100 3
16 74 473 282
7 5.000 V
7 5.000 V
3 GND
16 74 473 282
176160770 0
0
0
0
0
0
0
8
7 Pulser~
4 59 130 0 9 9
0 9 10 2 11 0 0 5 5 5
0
0 0 20528 0
0
2 V1
-7 -38 7 -30
0
0
0
0
0
0
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
8953 0 0
0
0
14 Logic Display~
6 382 23 0 1 3
11 8
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L1
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4441 0 0
0
0
14 Logic Display~
6 351 23 0 1 3
15 7
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L2
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3618 0 0
0
0
14 Logic Display~
6 321 23 0 1 3
14 6
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L3
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
14 Logic Display~
6 291 23 0 1 3
13 5
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L4
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5394 0 0
0
0
14 Logic Display~
6 261 23 0 1 3
12 4
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L5
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7734 0 0
0
0
14 Logic Display~
6 232 23 0 1 3
10 3
0
0 0 53344 0
6 100MEG
3 -16 45 -8
2 L6
17 -26 31 -18
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
9 Data Seq~
170 151 94 0 17 21
0 12 13 3 4 5 6 7 8 2
14 6 1 10 1 1 1 11
0
0 0 4208 0
6 DIGSRC
-21 -44 21 -36
3 DS1
-11 -54 10 -46
0
0
49 %D [%9i %10i][%1o %2o %3o %4o %5o %6o %7o %8o] %M
0
11 type:source
0
21

0 1 2 3 4 5 6 7 8 9
10 1 2 3 4 5 6 7 8 9
10 0
65 0 0 512 1 0 0 0
2 DS
3747 0 0
0
0
AAABACAEAIBACABAAIAEAC
7
9 3 2 0 0 4224 0 8 1 0 0 2
119 121
83 121
1 3 3 0 0 8320 0 7 8 0 0 3
232 41
232 85
183 85
4 1 4 0 0 4224 0 8 6 0 0 3
183 94
261 94
261 41
1 5 5 0 0 8320 0 5 8 0 0 3
291 41
291 103
183 103
6 1 6 0 0 4224 0 8 4 0 0 3
183 112
321 112
321 41
1 7 7 0 0 8320 0 3 8 0 0 3
351 41
351 121
183 121
8 1 8 0 0 4224 0 8 2 0 0 3
183 130
382 130
382 41
0
0
17 0 0
0
0
3 Vin
-1.5 -0.7 0.01
3 Vcc
10 14 1
100 0 1 100000
0 0.0005 2.5e-006 2.5e-006 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 100 100 0 0
98 66 608 126
0 0 0 0
608 66
98 66
608 66
608 126
0 0
1.01 0 0.495 0.009 1.01 1.01
12409 0
0 0.3 10
0
0 0 100 100 0 0
98 66 294 126
0 0 0 0
294 66
98 66
294 66
294 126
0 0
1e+007 1 12.16 12.184 1e+007 1e+007
12403 0
0 3e+006 5e+006
0
0 0 100 100 0 0
77 66 287 126
0 0 0 0
287 66
77 66
287 66
287 126
0 0
2000 1 2.38857 0 1999 1999
16 0
0 500 1000
0
0 0 100 100 0 0
98 66 296 126
0 0 0 0
296 66
98 66
296 66
296 126
0 0
1e+006 1 -3.55271e-015 0 999999 999999
12403 0
0 300000 500000
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0

CircuitMaker Text
5.5
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+009 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 20 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 9
0 71 1536 816
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
80 C:\Users\jonat\AppData\Local\Temp\Rar$EXa47972.16692\CIRCUIT MAKER_CM60S\BOM.DAT
0 7
0 71 1536 816
143654930 0
0
6 Title:
5 Name:
0
0
0
12
13 Logic Switch~
5 141 62 0 1 11
0 4
0
0 0 21344 270
2 0V
-6 -21 8 -13
1 C
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8953 0 0
0
0
13 Logic Switch~
5 115 57 0 1 11
0 3
0
0 0 21344 270
2 0V
-6 -21 8 -13
1 B
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4441 0 0
0
0
13 Logic Switch~
5 91 58 0 1 11
0 5
0
0 0 21344 270
2 0V
-6 -21 8 -13
1 A
-3 -31 4 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3618 0 0
0
0
14 Logic Display~
6 343 272 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6153 0 0
0
0
9 2-In XOR~
219 203 269 0 3 22
0 5 3 6
0
0 0 608 0
6 74LS86
-21 -24 21 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 6 0
1 U
5394 0 0
0
0
10 2-In XNOR~
219 281 301 0 3 22
0 6 4 2
0
0 0 608 0
4 4077
-7 -24 21 -16
3 U5A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
7734 0 0
0
0
14 Logic Display~
6 385 165 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9914 0 0
0
0
8 2-In OR~
219 240 174 0 3 22
0 5 3 8
0
0 0 608 0
6 74LS32
-21 -24 21 -16
3 U4A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3747 0 0
0
0
9 2-In NOR~
219 327 185 0 3 22
0 8 4 7
0
0 0 608 0
6 74LS02
-21 -24 21 -16
3 U3B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 3 2 1 5 6 4
8 9 10 11 12 13 0 0 0 0
0 6 0
65 0 0 0 4 2 3 0
1 U
3549 0 0
0
0
9 2-In AND~
219 251 101 0 3 22
0 5 3 10
0
0 0 608 0
6 74LS08
-21 -24 21 -16
3 U2A
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 2 0
1 U
7931 0 0
0
0
14 Logic Display~
6 372 87 0 1 2
10 9
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9325 0 0
0
0
10 2-In NAND~
219 315 110 0 3 22
0 10 4 9
0
0 0 608 0
6 74LS00
-14 -24 28 -16
3 U1B
-12 -25 9 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 4 5 6 1 2 3 4 5 6
10 9 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 2 1 0
1 U
8903 0 0
0
0
18
3 1 2 0 0 8320 0 6 4 0 0 3
320 301
343 301
343 290
0 2 3 0 0 4096 0 0 5 17 0 4
115 276
186 276
186 278
187 278
0 2 4 0 0 12288 0 0 6 16 0 4
141 307
172 307
172 310
265 310
0 1 5 0 0 4112 0 0 5 18 0 2
91 260
187 260
1 3 6 0 0 8320 0 6 5 0 0 3
265 292
265 269
236 269
1 3 7 0 0 8320 0 7 9 0 0 3
385 183
385 185
366 185
0 2 4 0 0 4096 0 0 9 16 0 4
141 199
278 199
278 194
314 194
1 3 8 0 0 4224 0 9 8 0 0 4
314 176
271 176
271 174
273 174
0 2 3 0 0 4096 0 0 8 17 0 4
115 182
202 182
202 183
227 183
0 1 5 0 0 4096 0 0 8 18 0 4
91 163
213 163
213 165
227 165
1 3 9 0 0 8320 0 11 12 0 0 3
372 105
372 110
342 110
3 1 10 0 0 4224 0 10 12 0 0 2
272 101
291 101
0 2 4 0 0 4096 0 0 12 16 0 3
141 127
291 127
291 119
0 2 3 0 0 4096 0 0 10 17 0 2
115 110
227 110
0 1 5 0 0 8192 0 0 10 18 0 3
91 89
91 92
227 92
1 0 4 0 0 4224 0 1 0 0 0 2
141 74
141 400
1 0 3 0 0 4224 0 2 0 0 0 2
115 69
115 399
1 0 5 0 0 4224 0 3 0 0 0 2
91 70
91 402
0
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
